module breadboard	();  

  

endmodule                           


module testbench();

  // Main code goes here
  
endmodule 































//Dr. Becker's cheat sheet of what is wrong in the code.
//The loop control variable can never reach 16, it is only 4 bits. Add another bit
//There needs to be a time dealy, such a #5, inside the for loop
