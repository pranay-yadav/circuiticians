/*
	Circuiticians Project Part 2
	CS 4341.001 Fall 2021 - University of Texas at Dallas
	
	Authors: 
		Jacob Medel, Christopher Clark, Donavin Sip, Pranay Yadav, Carlos Moran, Antonio Ramaj
	
*/



// Half Adder
module HalfAdder(a, b, carry, sum);

endmodule


// Full Adder
module FullAdder(a, b, carry, sum);
	
endmodule

// Adder-Subtracter
module AddSub(IN1, IN2, OP, S, CAR, OVF);

endmodule

// Multiplication
module Mul(IN1, IN2, P);

endmodule

// Division
module Div(IN1, IN2, Q, DE);

endmodule

// Modulo
module Mod(IN1, IN2, R, ME)

endmodule

// Decoder
module Dec(OP, SEL);

endmodule

// Multiplexer
module Mux(channels, SEL, OUT);

endmodule


module BreadBoard(IN1, IN2, OP, OUT, ERR);

endmodule


module TestBench();
 
endmodule  